module instruction_processor (clk,opcode,read_address1,read_address2,write_address,write_data,valid_address,read_data1,read_data2,done);
    input clk;
    input [2:0] opcode;
    output reg done;

    

    always @(posedge clk) begin
        
    end
endmodule